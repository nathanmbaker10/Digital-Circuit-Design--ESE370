*** SPICE deck for cell MemoryCellTest{sch} from library ESE370
*** Created on Fri Nov 19, 2021 15:30:10
*** Last revised on Sun Nov 21, 2021 20:44:10
*** Written on Sun Nov 21, 2021 20:44:19 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF
* Model cards are described in this file:
.include '~/Desktop/Shared VM (Desktop)/ESE370/22nm_HP.pm'

*** SUBCIRCUIT ESE370__inverter FROM CELL inverter{sch}
.SUBCKT ESE370__inverter a not_a_
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 not_a_ a gnd gnd N L=0.022U W=0.022U
Mpmos@0 vdd a not_a_ vdd P L=0.022U W=0.022U
.ENDS ESE370__inverter

*** SUBCIRCUIT ESE370__buffer FROM CELL buffer{sch}
.SUBCKT ESE370__buffer a out
** GLOBAL gnd
** GLOBAL vdd
Xinverter@0 a net@1 ESE370__inverter
Xinverter@1 net@1 out ESE370__inverter
.ENDS ESE370__buffer

*** SUBCIRCUIT ESE370__ColumnChooser FROM CELL ColumnChooser{sch}
.SUBCKT ESE370__ColumnChooser C0 C1 In
** GLOBAL gnd
** GLOBAL vdd
Xbuffer@0 In C1 ESE370__buffer
Xinverter@0 In C0 ESE370__inverter
.ENDS ESE370__ColumnChooser

*** SUBCIRCUIT ESE370__tri-state-buffer FROM CELL tri-state-buffer{sch}
.SUBCKT ESE370__tri-state-buffer En In out
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 out En net@24 gnd N L=0.022U W=0.022U
Mnmos@1 net@24 net@3 gnd gnd N L=0.022U W=0.022U
Mpmos@0 net@1 net@14 out vdd P L=0.022U W=0.022U
Mpmos@1 vdd net@3 net@1 vdd P L=0.022U W=0.022U
Xinverter@1 In net@3 ESE370__inverter
Xinverter@2 En net@14 ESE370__inverter
.ENDS ESE370__tri-state-buffer

*** SUBCIRCUIT ESE370__tristate-buffer-enable-inverted FROM CELL tristate-buffer-enable-inverted{sch}
.SUBCKT ESE370__tristate-buffer-enable-inverted en in out
** GLOBAL gnd
** GLOBAL vdd
Xinverter@0 en net@2 ESE370__inverter
Xtri-stat@0 net@2 in out ESE370__tri-state-buffer
.ENDS ESE370__tristate-buffer-enable-inverted

*** SUBCIRCUIT ESE370__ColumnDriver FROM CELL ColumnDriver{sch}
.SUBCKT ESE370__ColumnDriver b C D R/_Wr
** GLOBAL gnd
** GLOBAL vdd
Xtri-stat@0 C D net@25 ESE370__tri-state-buffer
Xtri-stat@1 C net@34 D ESE370__tri-state-buffer
Xtri-stat@2 R/_Wr net@25 b ESE370__tri-state-buffer
Xtristate@0 R/_Wr b net@34 ESE370__tristate-buffer-enable-inverted
.ENDS ESE370__ColumnDriver

*** SUBCIRCUIT ESE370__RAM_Cell FROM CELL RAM_Cell{sch}
.SUBCKT ESE370__RAM_Cell BL BL_ WL
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 net@0 WL BL gnd N L=0.022U W=0.022U
Mnmos@1 BL_ WL net@5 gnd N L=0.022U W=0.022U
Xinverter@0 net@0 net@5 ESE370__inverter
Xinverter@1 net@5 net@0 ESE370__inverter
.ENDS ESE370__RAM_Cell

*** SUBCIRCUIT ESE370__bitLineConditioning FROM CELL bitLineConditioning{sch}
.SUBCKT ESE370__bitLineConditioning BL BL_ CLK
** GLOBAL vdd
Mpmos@0 vdd CLK BL_ vdd P L=0.022U W=0.022U
Mpmos@1 BL CLK vdd vdd P L=0.022U W=0.022U
.ENDS ESE370__bitLineConditioning

*** SUBCIRCUIT ESE370__tristate-inverter FROM CELL tristate-inverter{sch}
.SUBCKT ESE370__tristate-inverter En In out
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 out In net@13 gnd N L=0.022U W=0.022U
Mnmos@1 net@13 En gnd gnd N L=0.022U W=0.022U
Mpmos@0 net@0 In out vdd P L=0.022U W=0.022U
Mpmos@1 vdd net@28 net@0 vdd P L=0.022U W=0.022U
Xinverter@2 En net@28 ESE370__inverter
.ENDS ESE370__tristate-inverter

*** SUBCIRCUIT ESE370__MemoryCellTester FROM CELL MemoryCellTester{sch}
.SUBCKT ESE370__MemoryCellTester PC Q Q_ Rd/Wr_ WL
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 net@39 WL vdd gnd N L=0.022U W=0.022U
XColumnCh@0 net@15 ColumnCh@0_C1 gnd ESE370__ColumnChooser
XColumnDr@0 net@12 net@15 Q Rd/Wr_ ESE370__ColumnDriver
XColumnDr@1 net@33 net@15 Q_ Rd/Wr_ ESE370__ColumnDriver
XRAM_Cell@0 net@12 net@33 net@39 ESE370__RAM_Cell
XbitLineC@0 net@12 net@33 net@79 ESE370__bitLineConditioning
Xtristate@0 Rd/Wr_ PC net@79 ESE370__tristate-inverter
.ENDS ESE370__MemoryCellTester

.global gnd vdd

*** TOP LEVEL CELL: MemoryCellTest{sch}
XMemoryCe@2 PC Q Q_ RW WL ESE370__MemoryCellTester
VVPWL@1 net@88 gnd pwl (0ns 0V) DC '0V' AC '0V' 0
VVPulse@2 PC gnd pulse (0 0.8V 0ns 10ps 10ps 33ps 333ps) DC '0V' AC '0V' 0
VVPulse@3 WL gnd pulse (0 0.8V 50ps 10ps 10ps 151.5ps 333ps) DC '0V' AC '0V' 0
VVPulse@4 RW gnd pulse (0 0.8V 333ps 10ps 10ps 666ps 1ns) DC '0V' AC '0V' 0
VV_Generi@0 vdd gnd DC 0.8 AC 0
Xinverter@4 net@88 net@99 ESE370__inverter
Xtristate@0 RW net@99 Q_ ESE370__tristate-buffer-enable-inverted
Xtristate@1 RW net@88 Q ESE370__tristate-buffer-enable-inverted
.END
