*** SPICE deck for cell nand2FO4{sch} from library ESE370
*** Created on Wed Sep 15, 2021 21:37:32
*** Last revised on Wed Sep 15, 2021 21:53:33
*** Written on Wed Sep 15, 2021 21:54:33 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF
* Model cards are described in this file:
.include '~/Desktop/Shared VM (Desktop)/ESE370/22nm_HP.pm'

*** SUBCIRCUIT ESE370__nand2 FROM CELL nand2{sch}
.SUBCKT ESE370__nand2 A B O
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 O A net@10 gnd N L=0.044U W=0.044U
Mnmos@1 net@10 B gnd gnd N L=0.044U W=0.044U
Mpmos@0 vdd A O vdd P L=0.044U W=0.044U
Mpmos@1 vdd B O vdd P L=0.044U W=0.044U
.ENDS ESE370__nand2

.global gnd vdd

*** TOP LEVEL CELL: nand2FO4{sch}
VVPulse@0 net@4 gnd pulse (0 0.8V 50ps 10ps 10ps 250ps 500ps) DC '0V' AC '0V' 0
VV_Generi@0 vdd gnd DC 0.8 AC 0
VV_Generi@1 net@7 gnd DC 0.8 AC 0
VV_Generi@2 net@16 gnd DC 0.8 AC 0
Xnand2@0 net@4 net@7 net@20 ESE370__nand2
Xnand2@1 net@20 net@16 nand2@1_O ESE370__nand2
Xnand2@2 net@20 net@16 net@37 ESE370__nand2
Xnand2@3 net@20 net@20 nand2@3_O ESE370__nand2
Xnand2@4 net@39 net@39 nand2@4_O ESE370__nand2
Xnand2@5 net@37 net@39 nand2@5_O ESE370__nand2
.END
