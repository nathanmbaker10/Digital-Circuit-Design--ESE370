*** SPICE deck for cell MemoryCellTesterInside{sch} from library ESE370
*** Created on Fri Nov 19, 2021 13:43:25
*** Last revised on Mon Nov 22, 2021 20:48:14
*** Written on Mon Nov 22, 2021 20:48:25 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF
* Model cards are described in this file:
.include C:\Users\shane\Downloads\22nm_HP.pm

*** SUBCIRCUIT ESE370__inverter FROM CELL inverter{sch}
.SUBCKT ESE370__inverter a not_a_
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 not_a_ a gnd gnd N L=0.022U W=0.022U
Mpmos@0 vdd a not_a_ vdd P L=0.022U W=0.022U
.ENDS ESE370__inverter

*** SUBCIRCUIT ESE370__tri-state-buffer FROM CELL tri-state-buffer{sch}
.SUBCKT ESE370__tri-state-buffer En In out
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 out En net@24 gnd N L=0.022U W=0.022U
Mnmos@1 net@24 net@3 gnd gnd N L=0.022U W=0.022U
Mpmos@0 net@1 net@14 out vdd P L=0.022U W=0.022U
Mpmos@1 vdd net@3 net@1 vdd P L=0.022U W=0.022U
Xinverter@1 In net@3 ESE370__inverter
Xinverter@2 En net@14 ESE370__inverter
.ENDS ESE370__tri-state-buffer

*** SUBCIRCUIT ESE370__tristate-buffer-enable-inverted FROM CELL tristate-buffer-enable-inverted{sch}
.SUBCKT ESE370__tristate-buffer-enable-inverted en in out
** GLOBAL gnd
** GLOBAL vdd
Xinverter@0 en net@2 ESE370__inverter
Xtri-stat@0 net@2 in out ESE370__tri-state-buffer
.ENDS ESE370__tristate-buffer-enable-inverted

*** SUBCIRCUIT ESE370__ColumnDriver FROM CELL ColumnDriver{sch}
.SUBCKT ESE370__ColumnDriver b d WR/_R
** GLOBAL gnd
** GLOBAL vdd
Xtri-stat@2 WR/_R d b ESE370__tri-state-buffer
Xtristate@0 WR/_R b d ESE370__tristate-buffer-enable-inverted
.ENDS ESE370__ColumnDriver

*** SUBCIRCUIT ESE370__RAM_Cell FROM CELL RAM_Cell{sch}
.SUBCKT ESE370__RAM_Cell BL BL_ WL
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 net@0 WL BL gnd N L=0.022U W=0.022U
Mnmos@1 BL_ WL net@5 gnd N L=0.022U W=0.022U
Xinverter@0 net@0 net@5 ESE370__inverter
Xinverter@1 net@5 net@0 ESE370__inverter
.ENDS ESE370__RAM_Cell

*** SUBCIRCUIT ESE370__bitLineConditioning FROM CELL bitLineConditioning{sch}
.SUBCKT ESE370__bitLineConditioning BL BL_ CLK
** GLOBAL vdd
Mpmos@0 vdd CLK BL_ vdd P L=0.022U W=0.022U
Mpmos@2 vdd CLK BL vdd P L=0.022U W=0.022U
.ENDS ESE370__bitLineConditioning

*** SUBCIRCUIT ESE370__tristate-inverter FROM CELL tristate-inverter{sch}
.SUBCKT ESE370__tristate-inverter En In out
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 out In net@13 gnd N L=0.022U W=0.022U
Mnmos@1 net@13 En gnd gnd N L=0.022U W=0.022U
Mpmos@0 net@0 In out vdd P L=0.022U W=0.022U
Mpmos@1 vdd net@28 net@0 vdd P L=0.022U W=0.022U
Xinverter@2 En net@28 ESE370__inverter
.ENDS ESE370__tristate-inverter

.global gnd vdd

*** TOP LEVEL CELL: MemoryCellTesterInside{sch}
XColumnDr@4 BL Q vdd ESE370__ColumnDriver
XColumnDr@5 BL_ Q_ vdd ESE370__ColumnDriver
XRAM_Cell@0 BL BL_ WL ESE370__RAM_Cell
VVPWL@0 net@365 gnd pwl (0ns 0.8 333ps 0.8 333ps 0 1ns 0 1ns 0.8 166ps 0.8) DC 0V AC 0V 0
VVPulse@1 PC gnd pulse (0.8V 0V 20ps 10ps 10ps 80ps 333ps) DC 0V AC 0V 0
VVPulse@2 net@380 gnd pulse (0V 0.8V 0ps 10ps 10ps 333ps 1ns) DC 0V AC 0V 0
VVPulse@3 WL gnd pulse (0 0.8V 50ps 10ps 10ps 151.5ps 333ps) DC 0V AC 0V 0
VV_Generi@0 vdd gnd DC 0.8 AC 0
XbitLineC@0 net@233 net@235 PC ESE370__bitLineConditioning
Xtri-stat@0 vdd net@365 Q ESE370__tri-state-buffer
Xtristate@2 vdd net@235 BL_ ESE370__tristate-buffer-enable-inverted
Xtristate@3 vdd net@233 BL ESE370__tristate-buffer-enable-inverted
Xtristate@4 vdd net@365 Q_ ESE370__tristate-inverter
.END
