*** SPICE deck for cell RowDecoder{sch} from library ESE370
*** Created on Sun Nov 28, 2021 23:37:44
*** Last revised on Mon Nov 29, 2021 16:23:49
*** Written on Mon Nov 29, 2021 16:24:09 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF
* Model cards are described in this file:
.include C:\Users\shane\Downloads\22nm_HP.pm

*** SUBCIRCUIT ESE370__inverter FROM CELL inverter{sch}
.SUBCKT ESE370__inverter a not_a_
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 not_a_ a gnd gnd N L=0.022U W=0.022U
Mpmos@0 vdd a not_a_ vdd P L=0.022U W=0.022U
.ENDS ESE370__inverter

*** SUBCIRCUIT ESE370__nand2 FROM CELL nand2{sch}
.SUBCKT ESE370__nand2 A B O
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 O A net@10 gnd N L=0.022U W=0.022U
Mnmos@1 net@10 B gnd gnd N L=0.022U W=0.022U
Mpmos@0 vdd A O vdd P L=0.022U W=0.022U
Mpmos@1 vdd B O vdd P L=0.022U W=0.022U
.ENDS ESE370__nand2

*** SUBCIRCUIT ESE370__and2 FROM CELL and2{sch}
.SUBCKT ESE370__and2 a b output
** GLOBAL gnd
** GLOBAL vdd
Xinverter@0 net@25 output ESE370__inverter
Xnand2@0 a b net@25 ESE370__nand2
.ENDS ESE370__and2

.global gnd vdd

*** TOP LEVEL CELL: RowDecoder{sch}
Mnmos@0 net@346 net@33 gnd gnd N L=0.022U W=0.022U
Mnmos@2 net@267 net@33 gnd gnd N L=0.022U W=0.022U
Mnmos@3 net@49 net@51 gnd gnd N L=0.022U W=0.022U
Mnmos@7 net@269 net@51 gnd gnd N L=0.022U W=0.022U
Mnmos@8 net@70 net@72 gnd gnd N L=0.022U W=0.022U
Mnmos@11 net@81 net@72 gnd gnd N L=0.022U W=0.022U
Mnmos@12 net@85 net@97 gnd gnd N L=0.022U W=0.022U
Mnmos@15 net@341 net@97 gnd gnd N L=0.022U W=0.022U
Mnmos@16 net@125 net@281 net@346 gnd N L=0.022U W=0.022U
Mnmos@17 net@130 A0 net@267 gnd N L=0.022U W=0.022U
Mnmos@18 net@139 net@281 net@49 gnd N L=0.022U W=0.022U
Mnmos@19 net@145 A0 net@269 gnd N L=0.022U W=0.022U
Mnmos@20 net@149 net@281 net@70 gnd N L=0.022U W=0.022U
Mnmos@21 net@153 A0 net@81 gnd N L=0.022U W=0.022U
Mnmos@22 net@161 net@281 net@85 gnd N L=0.022U W=0.022U
Mnmos@23 net@94 A0 net@341 gnd N L=0.022U W=0.022U
Mpmos@8 vdd net@208 net@125 vdd P L=0.022U W=0.022U
Mpmos@9 vdd net@208 net@130 vdd P L=0.022U W=0.022U
Mpmos@10 vdd net@208 net@139 vdd P L=0.022U W=0.022U
Mpmos@11 vdd net@208 net@145 vdd P L=0.022U W=0.022U
Mpmos@12 vdd net@208 net@149 vdd P L=0.022U W=0.022U
Mpmos@13 vdd net@208 net@153 vdd P L=0.022U W=0.022U
Mpmos@14 vdd net@208 net@161 vdd P L=0.022U W=0.022U
Mpmos@15 vdd net@208 net@94 vdd P L=0.022U W=0.022U
VVPulse@0 net@208 gnd pulse (0.8 0V 0ns 10ps 10ps 150ps 500ps) DC 0V AC 0V 0
VVPulse@1 A0 gnd pulse (0.8 0V 0ps 10ps 10ps 500ps 1000ps) DC 0V AC 0V 0
VVPulse@2 A1 gnd pulse (0.8 0V 0ps 10ps 10ps 1000ps 2000ps) DC 0V AC 0V 0
VVPulse@3 A2 gnd pulse (0.8 0V 0ps 10ps 10ps 2000ps 4000ps) DC 0V AC 0V 0
VV_Generi@0 vdd gnd DC 0.8 AC 0
Xand2@0 A2 A1 net@97 ESE370__and2
Xand2@1 net@10 A1 net@51 ESE370__and2
Xand2@2 A2 net@9 net@72 ESE370__and2
Xand2@3 net@8 net@7 net@33 ESE370__and2
Xinverter@1 A1 net@7 ESE370__inverter
Xinverter@2 A2 net@8 ESE370__inverter
Xinverter@3 A1 net@9 ESE370__inverter
Xinverter@4 A2 net@10 ESE370__inverter
Xinverter@6 net@125 WL0 ESE370__inverter
Xinverter@7 net@130 WL1 ESE370__inverter
Xinverter@8 net@139 WL2 ESE370__inverter
Xinverter@9 net@145 WL3 ESE370__inverter
Xinverter@10 net@149 WL4 ESE370__inverter
Xinverter@11 net@153 WL5 ESE370__inverter
Xinverter@12 net@161 WL6 ESE370__inverter
Xinverter@13 net@94 WL7 ESE370__inverter
Xinverter@14 A0 net@281 ESE370__inverter
.END
