*** SPICE deck for cell SRAMtests{sch} from library ESE370
*** Created on Thu Dec 02, 2021 20:42:33
*** Last revised on Fri Dec 03, 2021 00:37:49
*** Written on Fri Dec 03, 2021 02:04:24 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF
* Model cards are described in this file:
.include '~/Desktop/Shared VM (Desktop)/ESE370/22nm_HP.pm'

*** SUBCIRCUIT ESE370__inverter FROM CELL inverter{sch}
.SUBCKT ESE370__inverter a not_a_
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 not_a_ a gnd gnd N L=0.022U W=0.022U
Mpmos@0 vdd a not_a_ vdd P L=0.022U W=0.022U
.ENDS ESE370__inverter

*** SUBCIRCUIT ESE370__buffer FROM CELL buffer{sch}
.SUBCKT ESE370__buffer a out
** GLOBAL gnd
** GLOBAL vdd
Xinverter@0 a net@1 ESE370__inverter
Xinverter@1 net@1 out ESE370__inverter
.ENDS ESE370__buffer

*** SUBCIRCUIT ESE370__ColumnChooser FROM CELL ColumnChooser{sch}
.SUBCKT ESE370__ColumnChooser C0 C1 In
** GLOBAL gnd
** GLOBAL vdd
Xbuffer@0 In C1 ESE370__buffer
Xinverter@0 In C0 ESE370__inverter
.ENDS ESE370__ColumnChooser

*** SUBCIRCUIT ESE370__tri-state-buffer FROM CELL tri-state-buffer{sch}
.SUBCKT ESE370__tri-state-buffer En In out
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 out En net@24 gnd N L=0.022U W=0.022U
Mnmos@1 net@24 net@3 gnd gnd N L=0.022U W=0.022U
Mpmos@0 net@1 net@14 out vdd P L=0.022U W=0.022U
Mpmos@1 vdd net@3 net@1 vdd P L=0.022U W=0.022U
Xinverter@1 In net@3 ESE370__inverter
Xinverter@2 En net@14 ESE370__inverter
.ENDS ESE370__tri-state-buffer

*** SUBCIRCUIT ESE370__tristate-buffer-enable-inverted FROM CELL tristate-buffer-enable-inverted{sch}
.SUBCKT ESE370__tristate-buffer-enable-inverted en in out
** GLOBAL gnd
** GLOBAL vdd
Xinverter@0 en net@2 ESE370__inverter
Xtri-stat@0 net@2 in out ESE370__tri-state-buffer
.ENDS ESE370__tristate-buffer-enable-inverted

*** SUBCIRCUIT ESE370__ColumnDriver FROM CELL ColumnDriver{sch}
.SUBCKT ESE370__ColumnDriver b Cin d WR/_R
** GLOBAL gnd
** GLOBAL vdd
Xtri-stat@0 WR/_R d net@162 ESE370__tri-state-buffer
Xtri-stat@1 Cin net@162 b ESE370__tri-state-buffer
Xtri-stat@2 Cin b net@181 ESE370__tri-state-buffer
Xtristate@8 WR/_R net@181 net@187 ESE370__tristate-buffer-enable-inverted
.ENDS ESE370__ColumnDriver

*** SUBCIRCUIT ESE370__ColumnDecoderBus FROM CELL ColumnDecoderBus{sch}
.SUBCKT ESE370__ColumnDecoderBus BL_[7] BL_[6] BL_[5] BL_[4] BL_[3] BL_[2] BL_[1] BL_[0] BL[7] BL[6] BL[5] BL[4] BL[3] BL[2] BL[1] BL[0] Cin D_[3] D_[2] D_[1] D_[0] D[3] D[2] D[1] D[0] Wr/_R
** GLOBAL gnd
** GLOBAL vdd
XColumnCh@0 net@8 net@46 Cin ESE370__ColumnChooser
XColumnDr@0 BL[0] net@8 D[0] Wr/_R ESE370__ColumnDriver
XColumnDr@1 BL_[0] net@8 D_[0] Wr/_R ESE370__ColumnDriver
XColumnDr@4 BL[1] net@8 D[1] Wr/_R ESE370__ColumnDriver
XColumnDr@5 BL_[1] net@8 D_[1] Wr/_R ESE370__ColumnDriver
XColumnDr@6 BL[2] net@8 D[2] Wr/_R ESE370__ColumnDriver
XColumnDr@7 BL_[2] net@8 D_[2] Wr/_R ESE370__ColumnDriver
XColumnDr@8 BL[3] net@8 D[3] Wr/_R ESE370__ColumnDriver
XColumnDr@9 BL_[3] net@8 D_[3] Wr/_R ESE370__ColumnDriver
XColumnDr@10 BL[4] net@46 D[0] Wr/_R ESE370__ColumnDriver
XColumnDr@11 BL_[4] net@46 D_[0] Wr/_R ESE370__ColumnDriver
XColumnDr@12 BL[5] net@46 D[1] Wr/_R ESE370__ColumnDriver
XColumnDr@13 BL_[5] net@46 D_[1] Wr/_R ESE370__ColumnDriver
XColumnDr@14 BL[6] net@46 D[2] Wr/_R ESE370__ColumnDriver
XColumnDr@15 BL_[6] net@46 D_[2] Wr/_R ESE370__ColumnDriver
XColumnDr@16 BL[7] net@46 D[3] Wr/_R ESE370__ColumnDriver
XColumnDr@17 BL_[7] net@46 D_[3] Wr/_R ESE370__ColumnDriver
.ENDS ESE370__ColumnDecoderBus

*** SUBCIRCUIT ESE370__RAM_Cell FROM CELL RAM_Cell{sch}
.SUBCKT ESE370__RAM_Cell BL BL_ WL
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 net@0 WL BL gnd N L=0.022U W=0.044U
Mnmos@1 BL_ WL net@10 gnd N L=0.022U W=0.022U
Mnmos@2 net@10 net@0 gnd gnd N L=0.022U W=0.044U
Mnmos@3 net@0 net@10 gnd gnd N L=0.022U W=0.022U
Mpmos@0 vdd net@0 net@10 vdd P L=0.022U W=0.022U
Mpmos@1 vdd net@10 net@0 vdd P L=0.022U W=0.022U
.ENDS ESE370__RAM_Cell

*** SUBCIRCUIT ESE370__nand2 FROM CELL nand2{sch}
.SUBCKT ESE370__nand2 A B O
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 O A net@10 gnd N L=0.022U W=0.022U
Mnmos@1 net@10 B gnd gnd N L=0.022U W=0.022U
Mpmos@0 vdd A O vdd P L=0.022U W=0.022U
Mpmos@1 vdd B O vdd P L=0.022U W=0.022U
.ENDS ESE370__nand2

*** SUBCIRCUIT ESE370__and2 FROM CELL and2{sch}
.SUBCKT ESE370__and2 a b output
** GLOBAL gnd
** GLOBAL vdd
Xinverter@0 net@25 output ESE370__inverter
Xnand2@0 a b net@25 ESE370__nand2
.ENDS ESE370__and2

*** SUBCIRCUIT ESE370__RowDecoder FROM CELL RowDecoder{sch}
.SUBCKT ESE370__RowDecoder Addr[2] Addr[1] Addr[0] WL0 WL1 WL2 WL3 WL4 WL5 WL6 WL7 _PC
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 net@346 net@33 gnd gnd N L=0.022U W=0.022U
Mnmos@2 net@267 net@33 gnd gnd N L=0.022U W=0.022U
Mnmos@3 net@49 net@51 gnd gnd N L=0.022U W=0.022U
Mnmos@7 net@269 net@51 gnd gnd N L=0.022U W=0.022U
Mnmos@8 net@70 net@72 gnd gnd N L=0.022U W=0.022U
Mnmos@11 net@81 net@72 gnd gnd N L=0.022U W=0.022U
Mnmos@12 net@85 net@97 gnd gnd N L=0.022U W=0.022U
Mnmos@15 net@341 net@97 gnd gnd N L=0.022U W=0.022U
Mnmos@16 net@125 net@281 net@346 gnd N L=0.022U W=0.022U
Mnmos@17 net@130 Addr[0] net@267 gnd N L=0.022U W=0.022U
Mnmos@18 net@139 net@281 net@49 gnd N L=0.022U W=0.022U
Mnmos@19 net@145 Addr[0] net@269 gnd N L=0.022U W=0.022U
Mnmos@20 net@149 net@281 net@70 gnd N L=0.022U W=0.022U
Mnmos@21 net@153 Addr[0] net@81 gnd N L=0.022U W=0.022U
Mnmos@22 net@161 net@281 net@85 gnd N L=0.022U W=0.022U
Mnmos@23 net@94 Addr[0] net@341 gnd N L=0.022U W=0.022U
Mpmos@8 vdd _PC net@125 vdd P L=0.022U W=0.044U
Mpmos@9 vdd _PC net@130 vdd P L=0.022U W=0.044U
Mpmos@10 vdd _PC net@139 vdd P L=0.022U W=0.044U
Mpmos@11 vdd _PC net@145 vdd P L=0.022U W=0.044U
Mpmos@12 vdd _PC net@149 vdd P L=0.022U W=0.044U
Mpmos@13 vdd _PC net@153 vdd P L=0.022U W=0.044U
Mpmos@14 vdd _PC net@161 vdd P L=0.022U W=0.044U
Mpmos@15 vdd _PC net@94 vdd P L=0.022U W=0.044U
Xand2@0 Addr[1] Addr[2] net@97 ESE370__and2
Xand2@1 net@10 Addr[2] net@51 ESE370__and2
Xand2@2 Addr[1] net@9 net@72 ESE370__and2
Xand2@3 net@8 net@7 net@33 ESE370__and2
Xinverter@1 Addr[2] net@7 ESE370__inverter
Xinverter@2 Addr[1] net@8 ESE370__inverter
Xinverter@3 Addr[2] net@9 ESE370__inverter
Xinverter@4 Addr[1] net@10 ESE370__inverter
Xinverter@6 net@125 WL0 ESE370__inverter
Xinverter@7 net@130 WL1 ESE370__inverter
Xinverter@8 net@139 WL2 ESE370__inverter
Xinverter@9 net@145 WL3 ESE370__inverter
Xinverter@10 net@149 WL4 ESE370__inverter
Xinverter@11 net@153 WL5 ESE370__inverter
Xinverter@12 net@161 WL6 ESE370__inverter
Xinverter@13 net@94 WL7 ESE370__inverter
Xinverter@14 Addr[0] net@281 ESE370__inverter
.ENDS ESE370__RowDecoder

*** SUBCIRCUIT ESE370__bitLineConditioning FROM CELL bitLineConditioning{sch}
.SUBCKT ESE370__bitLineConditioning BL BL_ CLK
** GLOBAL vdd
Mpmos@0 vdd CLK BL_ vdd P L=0.022U W=0.022U
Mpmos@2 vdd CLK BL vdd P L=0.022U W=0.022U
.ENDS ESE370__bitLineConditioning

*** SUBCIRCUIT ESE370__SRAM FROM CELL SRAM{sch}
.SUBCKT ESE370__SRAM Addr[3] Addr[2] Addr[1] Addr[0] bl0 D_[3] D_[2] D_[1] D_[0] D[3] D[2] D[1] D[0] PC pcafter wl0 wl1 WR/_R
** GLOBAL gnd
** GLOBAL vdd
XColumnDe@0 net@161 net@147 net@133 net@119 bl_4 bl_3 bl_2 bl_ net@154 net@140 net@126 net@112 bl4 bl3 bl2 bl0 Addr[3] D_[0] D_[1] D_[2] D_[3] D[0] D[1] D[2] D[3] WR/_R ESE370__ColumnDecoderBus
XRAM_Cell@0 bl0 bl_ wl0 ESE370__RAM_Cell
XRAM_Cell@1 bl2 bl_2 wl0 ESE370__RAM_Cell
XRAM_Cell@2 bl3 bl_3 wl0 ESE370__RAM_Cell
XRAM_Cell@3 bl4 bl_4 wl0 ESE370__RAM_Cell
XRAM_Cell@8 net@112 net@119 wl0 ESE370__RAM_Cell
XRAM_Cell@9 net@126 net@133 wl0 ESE370__RAM_Cell
XRAM_Cell@10 net@140 net@147 wl0 ESE370__RAM_Cell
XRAM_Cell@11 net@154 net@161 wl0 ESE370__RAM_Cell
XRAM_Cell@12 bl0 bl_ wl1 ESE370__RAM_Cell
XRAM_Cell@13 bl2 bl_2 wl1 ESE370__RAM_Cell
XRAM_Cell@14 bl3 bl_3 wl1 ESE370__RAM_Cell
XRAM_Cell@15 bl4 bl_4 wl1 ESE370__RAM_Cell
XRAM_Cell@16 net@112 net@119 wl1 ESE370__RAM_Cell
XRAM_Cell@17 net@126 net@133 wl1 ESE370__RAM_Cell
XRAM_Cell@18 net@140 net@147 wl1 ESE370__RAM_Cell
XRAM_Cell@19 net@154 net@161 wl1 ESE370__RAM_Cell
XRAM_Cell@20 bl0 bl_ wl2 ESE370__RAM_Cell
XRAM_Cell@21 bl2 bl_2 wl2 ESE370__RAM_Cell
XRAM_Cell@22 bl3 bl_3 wl2 ESE370__RAM_Cell
XRAM_Cell@23 bl4 bl_4 wl2 ESE370__RAM_Cell
XRAM_Cell@24 net@112 net@119 wl2 ESE370__RAM_Cell
XRAM_Cell@25 net@126 net@133 wl2 ESE370__RAM_Cell
XRAM_Cell@26 net@140 net@147 wl2 ESE370__RAM_Cell
XRAM_Cell@27 net@154 net@161 wl2 ESE370__RAM_Cell
XRAM_Cell@28 bl0 bl_ wl3 ESE370__RAM_Cell
XRAM_Cell@29 bl2 bl_2 wl3 ESE370__RAM_Cell
XRAM_Cell@30 bl3 bl_3 wl3 ESE370__RAM_Cell
XRAM_Cell@31 bl4 bl_4 wl3 ESE370__RAM_Cell
XRAM_Cell@32 net@112 net@119 wl3 ESE370__RAM_Cell
XRAM_Cell@33 net@126 net@133 wl3 ESE370__RAM_Cell
XRAM_Cell@34 net@140 net@147 wl3 ESE370__RAM_Cell
XRAM_Cell@35 net@154 net@161 wl3 ESE370__RAM_Cell
XRAM_Cell@36 bl0 bl_ wl4 ESE370__RAM_Cell
XRAM_Cell@37 bl2 bl_2 wl4 ESE370__RAM_Cell
XRAM_Cell@38 bl3 bl_3 wl4 ESE370__RAM_Cell
XRAM_Cell@39 bl4 bl_4 wl4 ESE370__RAM_Cell
XRAM_Cell@40 net@112 net@119 wl4 ESE370__RAM_Cell
XRAM_Cell@41 net@126 net@133 wl4 ESE370__RAM_Cell
XRAM_Cell@42 net@140 net@147 wl4 ESE370__RAM_Cell
XRAM_Cell@43 net@154 net@161 wl4 ESE370__RAM_Cell
XRAM_Cell@44 bl0 bl_ wl5 ESE370__RAM_Cell
XRAM_Cell@45 bl2 bl_2 wl5 ESE370__RAM_Cell
XRAM_Cell@46 bl3 bl_3 wl5 ESE370__RAM_Cell
XRAM_Cell@47 bl4 bl_4 wl5 ESE370__RAM_Cell
XRAM_Cell@48 net@112 net@119 wl5 ESE370__RAM_Cell
XRAM_Cell@49 net@126 net@133 wl5 ESE370__RAM_Cell
XRAM_Cell@50 net@140 net@147 wl5 ESE370__RAM_Cell
XRAM_Cell@51 net@154 net@161 wl5 ESE370__RAM_Cell
XRAM_Cell@52 bl0 bl_ wl6 ESE370__RAM_Cell
XRAM_Cell@53 bl2 bl_2 wl6 ESE370__RAM_Cell
XRAM_Cell@54 bl3 bl_3 wl6 ESE370__RAM_Cell
XRAM_Cell@55 bl4 bl_4 wl6 ESE370__RAM_Cell
XRAM_Cell@56 net@112 net@119 wl6 ESE370__RAM_Cell
XRAM_Cell@57 net@126 net@133 wl6 ESE370__RAM_Cell
XRAM_Cell@58 net@140 net@147 wl6 ESE370__RAM_Cell
XRAM_Cell@59 net@154 net@161 wl6 ESE370__RAM_Cell
XRAM_Cell@60 bl0 bl_ wl7 ESE370__RAM_Cell
XRAM_Cell@61 bl2 bl_2 wl7 ESE370__RAM_Cell
XRAM_Cell@62 bl3 bl_3 wl7 ESE370__RAM_Cell
XRAM_Cell@63 bl4 bl_4 wl7 ESE370__RAM_Cell
XRAM_Cell@64 net@112 net@119 wl7 ESE370__RAM_Cell
XRAM_Cell@65 net@126 net@133 wl7 ESE370__RAM_Cell
XRAM_Cell@66 net@140 net@147 wl7 ESE370__RAM_Cell
XRAM_Cell@67 net@154 net@161 wl7 ESE370__RAM_Cell
XRowDecod@4 Addr[2] Addr[1] Addr[0] wl0 wl1 wl2 wl3 wl4 wl5 wl6 wl7 PC ESE370__RowDecoder
XbitLineC@0 bl0 bl_ pcafter ESE370__bitLineConditioning
XbitLineC@1 bl2 bl_2 pcafter ESE370__bitLineConditioning
XbitLineC@2 bl3 bl_3 pcafter ESE370__bitLineConditioning
XbitLineC@3 bl4 bl_4 pcafter ESE370__bitLineConditioning
XbitLineC@4 net@112 net@119 pcafter ESE370__bitLineConditioning
XbitLineC@5 net@126 net@133 pcafter ESE370__bitLineConditioning
XbitLineC@7 net@140 net@147 pcafter ESE370__bitLineConditioning
XbitLineC@8 net@154 net@161 pcafter ESE370__bitLineConditioning
Xtristate@1 WR/_R PC pcafter ESE370__tristate-buffer-enable-inverted
.ENDS ESE370__SRAM

*** SUBCIRCUIT ESE370__4buffers FROM CELL 4buffers{sch}
.SUBCKT ESE370__4buffers A B
** GLOBAL gnd
** GLOBAL vdd
Xbuffer@0 A net@0 ESE370__buffer
Xbuffer@1 net@0 net@1 ESE370__buffer
Xbuffer@2 net@1 net@2 ESE370__buffer
Xbuffer@3 net@2 B ESE370__buffer
.ENDS ESE370__4buffers

*** SUBCIRCUIT ESE370__AddressSelector FROM CELL AddressSelector{sch}
.SUBCKT ESE370__AddressSelector Addr0 Addr1 Addr2 Addr3 Raddr0 Raddr1 Raddr2 Raddr3 Wr/_RCtrl Wraddr0 Wraddr1 Wraddr2 Wraddr3
** GLOBAL gnd
** GLOBAL vdd
Xtri-stat@0 Wr/_RCtrl Wraddr0 Addr0 ESE370__tri-state-buffer
Xtri-stat@1 Wr/_RCtrl Wraddr1 Addr1 ESE370__tri-state-buffer
Xtri-stat@2 Wr/_RCtrl Wraddr2 Addr2 ESE370__tri-state-buffer
Xtri-stat@3 Wr/_RCtrl Wraddr3 Addr3 ESE370__tri-state-buffer
Xtristate@0 Wr/_RCtrl Raddr0 Addr0 ESE370__tristate-buffer-enable-inverted
Xtristate@1 Wr/_RCtrl Raddr1 Addr1 ESE370__tristate-buffer-enable-inverted
Xtristate@2 Wr/_RCtrl Raddr2 Addr2 ESE370__tristate-buffer-enable-inverted
Xtristate@3 Wr/_RCtrl Raddr3 Addr3 ESE370__tristate-buffer-enable-inverted
.ENDS ESE370__AddressSelector

*** SUBCIRCUIT ESE370__nor2 FROM CELL nor2{sch}
.SUBCKT ESE370__nor2 a b o
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 o b gnd gnd N L=0.022U W=0.022U
Mnmos@1 o a gnd gnd N L=0.022U W=0.022U
Mpmos@0 vdd a net@12 vdd P L=0.022U W=0.022U
Mpmos@1 net@12 b o vdd P L=0.022U W=0.022U
.ENDS ESE370__nor2

*** SUBCIRCUIT ESE370__2phaseclock FROM CELL 2phaseclock{sch}
.SUBCKT ESE370__2phaseclock clock1 clock2 in
** GLOBAL gnd
** GLOBAL vdd
Xbuffer@0 in net@5 ESE370__buffer
Xinverter@0 in net@4 ESE370__inverter
Xnor2@0 net@4 clock2 clock1 ESE370__nor2
Xnor2@1 clock1 net@5 clock2 ESE370__nor2
.ENDS ESE370__2phaseclock

*** SUBCIRCUIT ESE370__3nandlatch FROM CELL 3nandlatch{sch}
.SUBCKT ESE370__3nandlatch clock in out
** GLOBAL gnd
** GLOBAL vdd
Xinverter@0 clock net@6 ESE370__inverter
Xnand2@0 in clock net@8 ESE370__nand2
Xnand2@1 net@6 out net@10 ESE370__nand2
Xnand2@2 net@8 net@10 out ESE370__nand2
.ENDS ESE370__3nandlatch

*** SUBCIRCUIT ESE370__PositiveRegister FROM CELL PositiveRegister{sch}
.SUBCKT ESE370__PositiveRegister clk d q
** GLOBAL gnd
** GLOBAL vdd
X_2phasecl@0 net@20 net@24 clk ESE370__2phaseclock
X_3nandlat@0 net@24 d net@0 ESE370__3nandlatch
X_3nandlat@1 net@20 net@0 q ESE370__3nandlatch
.ENDS ESE370__PositiveRegister

*** SUBCIRCUIT ESE370__XNOR_PT FROM CELL XNOR_PT{sch}
.SUBCKT ESE370__XNOR_PT A B out
** GLOBAL gnd
** GLOBAL vdd
Mnmos@2 net@53 net@39 B gnd N L=0.022U W=0.022U
Mnmos@3 net@53 A net@44 gnd N L=0.022U W=0.022U
Xbuffer@0 net@58 out ESE370__buffer
Xinverter@0 A net@39 ESE370__inverter
Xinverter@1 B net@44 ESE370__inverter
Xinverter@2 net@53 net@58 ESE370__inverter
.ENDS ESE370__XNOR_PT

*** SUBCIRCUIT ESE370__inverter1 FROM CELL inverter1{sch}
.SUBCKT ESE370__inverter1 a not_a_
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 not_a_ a gnd gnd N L=0.022U W=0.198U
Mpmos@0 vdd a not_a_ vdd P L=0.022U W=0.614U
.ENDS ESE370__inverter1

*** SUBCIRCUIT ESE370__nand2_sized FROM CELL nand2_sized{sch}
.SUBCKT ESE370__nand2_sized A B O
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 O A net@10 gnd N L=0.022U W=0.022U
Mnmos@1 net@10 B gnd gnd N L=0.022U W=0.022U
Mpmos@0 vdd A O vdd P L=0.022U W=0.022U
Mpmos@1 vdd B O vdd P L=0.022U W=0.022U
.ENDS ESE370__nand2_sized

*** SUBCIRCUIT ESE370__and2_sized FROM CELL and2_sized{sch}
.SUBCKT ESE370__and2_sized a b output
** GLOBAL gnd
** GLOBAL vdd
Xinverter@2 net@45 output ESE370__inverter1
Xnand2_si@0 a b net@45 ESE370__nand2_sized
.ENDS ESE370__and2_sized

*** SUBCIRCUIT ESE370__Readaddr__Wraddr FROM CELL Readaddr==Wraddr{sch}
.SUBCKT ESE370__Readaddr__Wraddr Radd__WRadd rdAddr0 rdaddr1 rdaddr2 rdaddr3 wraddr0 wraddr1 wraddr2 wraddr3
** GLOBAL gnd
** GLOBAL vdd
XXNOR_PT@1 rdAddr0 wraddr0 net@0 ESE370__XNOR_PT
XXNOR_PT@2 rdaddr1 wraddr1 net@3 ESE370__XNOR_PT
XXNOR_PT@3 rdaddr2 wraddr2 net@5 ESE370__XNOR_PT
XXNOR_PT@4 rdaddr3 wraddr3 net@7 ESE370__XNOR_PT
Xand2@0 net@9 net@11 Radd__WRadd ESE370__and2
Xand2_siz@0 net@0 net@3 net@9 ESE370__and2_sized
Xand2_siz@1 net@5 net@7 net@11 ESE370__and2_sized
.ENDS ESE370__Readaddr__Wraddr

*** SUBCIRCUIT ESE370__TristateBufferSized FROM CELL TristateBufferSized{sch}
.SUBCKT ESE370__TristateBufferSized En In out
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 out En net@6 gnd N L=0.022U W=0.088U
Mnmos@1 net@6 net@10 gnd gnd N L=0.022U W=0.088U
Mpmos@0 net@1 net@17 out vdd P L=0.022U W=0.088U
Mpmos@1 vdd net@10 net@1 vdd P L=0.022U W=0.088U
Xinverter@0 In net@10 ESE370__inverter
Xinverter@1 En net@17 ESE370__inverter
.ENDS ESE370__TristateBufferSized

*** SUBCIRCUIT ESE370__4bitReg FROM CELL 4bitReg{sch}
.SUBCKT ESE370__4bitReg CLK In[3] In[2] In[1] In[0] Out[3] Out[2] Out[1] Out[0]
** GLOBAL gnd
** GLOBAL vdd
XPositive@1 CLK In[3] Out[3] ESE370__PositiveRegister
XPositive@2 CLK In[2] Out[2] ESE370__PositiveRegister
XPositive@3 CLK In[1] Out[1] ESE370__PositiveRegister
XPositive@4 CLK In[0] Out[0] ESE370__PositiveRegister
.ENDS ESE370__4bitReg

*** SUBCIRCUIT ESE370__NAND2sized FROM CELL NAND2sized{sch}
.SUBCKT ESE370__NAND2sized A B out
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 net@1 B gnd gnd N L=0.022U W=0.11U
Mnmos@1 out A net@1 gnd N L=0.022U W=0.11U
Mpmos@0 vdd A out vdd P L=0.022U W=0.176U
Mpmos@1 vdd B out vdd P L=0.022U W=0.176U
.ENDS ESE370__NAND2sized

*** SUBCIRCUIT ESE370__nand2dc FROM CELL nand2dc{sch}
.SUBCKT ESE370__nand2dc A B out
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 net@1 B gnd gnd N L=0.022U W=0.022U
Mnmos@1 out A net@1 gnd N L=0.022U W=0.022U
Mpmos@2 vdd A out vdd P L=0.022U W=0.022U
Mpmos@3 vdd B out vdd P L=0.022U W=0.022U
.ENDS ESE370__nand2dc

*** SUBCIRCUIT ESE370__newXOR FROM CELL newXOR{sch}
.SUBCKT ESE370__newXOR A B out
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 out A net@18 gnd N L=0.022U W=0.022U
Mnmos@1 out net@46 net@19 gnd N L=0.022U W=0.022U
Mnmos@2 net@18 B gnd gnd N L=0.022U W=0.022U
Mnmos@3 net@19 net@51 gnd gnd N L=0.022U W=0.022U
Mpmos@0 vdd net@46 net@8 vdd P L=0.022U W=0.022U
Mpmos@1 vdd A net@7 vdd P L=0.022U W=0.022U
Mpmos@2 net@8 B out vdd P L=0.022U W=0.022U
Mpmos@3 net@7 net@51 out vdd P L=0.022U W=0.022U
Xinverter@0 A net@46 ESE370__inverter
Xinverter@1 B net@51 ESE370__inverter
.ENDS ESE370__newXOR

*** SUBCIRCUIT ESE370__Standardadder FROM CELL Standardadder{sch}
.SUBCKT ESE370__Standardadder A B Cin Cout S
** GLOBAL gnd
** GLOBAL vdd
XNAND2siz@0 net@36 Cin net@51 ESE370__NAND2sized
XNAND2siz@1 net@51 net@53 Cout ESE370__NAND2sized
Xnand2dc@0 A B net@53 ESE370__nand2dc
XnewXOR@0 A B net@36 ESE370__newXOR
XnewXOR@1 net@36 Cin S ESE370__newXOR
.ENDS ESE370__Standardadder

*** SUBCIRCUIT ESE370__PlusOne FROM CELL PlusOne{sch}
.SUBCKT ESE370__PlusOne in0 in1 in2 in3 out0 out1 out2 out3
** GLOBAL gnd
** GLOBAL vdd
XStandard@0 in0 vdd gnd net@5 out0 ESE370__Standardadder
XStandard@1 in1 gnd net@5 net@6 out1 ESE370__Standardadder
XStandard@2 in2 gnd net@6 net@9 out2 ESE370__Standardadder
XStandard@3 in3 gnd net@9 Standard@3_Cout out3 ESE370__Standardadder
.ENDS ESE370__PlusOne

*** SUBCIRCUIT ESE370__addressLoop FROM CELL addressLoop{sch}
.SUBCKT ESE370__addressLoop Addr[3] Addr[2] Addr[1] Addr[0] clk En/Deq
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 net@6 pc gnd gnd N L=0.044U W=0.044U
Mnmos@1 net@3 pc gnd gnd N L=0.044U W=0.044U
Mnmos@2 net@38 pc gnd gnd N L=0.044U W=0.044U
Mnmos@3 net@1 pc gnd gnd N L=0.044U W=0.044U
X_4bitReg@0 clk net@1 net@38 net@3 net@6 Addr[3] Addr[2] Addr[1] Addr[0] ESE370__4bitReg
XPlusOne@0 Addr[0] Addr[1] Addr[2] Addr[3] net@18 net@20 net@24 net@25 ESE370__PlusOne
VVPulse@0 pc gnd pulse (0 0.8V 0ns 10ps 10ps 80ps 1s) DC '0V' AC '0V' 0
Xtri-stat@0 En/Deq net@20 net@3 ESE370__tri-state-buffer
Xtri-stat@1 En/Deq net@18 net@6 ESE370__tri-state-buffer
Xtri-stat@2 En/Deq net@24 net@38 ESE370__tri-state-buffer
Xtri-stat@3 En/Deq net@25 net@1 ESE370__tri-state-buffer
Xtristate@0 En/Deq Addr[3] net@1 ESE370__tristate-buffer-enable-inverted
Xtristate@1 En/Deq Addr[2] net@38 ESE370__tristate-buffer-enable-inverted
Xtristate@2 En/Deq Addr[1] net@3 ESE370__tristate-buffer-enable-inverted
Xtristate@3 En/Deq Addr[0] net@6 ESE370__tristate-buffer-enable-inverted
.ENDS ESE370__addressLoop

*** SUBCIRCUIT ESE370__controlLogic FROM CELL controlLogic{sch}
.SUBCKT ESE370__controlLogic Addr0 Addr1 Addr2 Addr3 clk DQ Empty_next ENQ Full_next WRCtrl
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 Last__write net@208 gnd gnd N L=0.044U W=0.044U
X_4buffers@2 net@287 net@309 ESE370__4buffers
XAddressS@0 Addr0 Addr1 Addr2 Addr3 rdaddr0 rdaddr1 rdaddr2 rdaddr3 net@309 wraddr0 wraddr1 wraddr2 wraddr3 ESE370__AddressSelector
XPositive@0 clk this__write Last__write ESE370__PositiveRegister
XReadaddr@0 ptrflag wraddr0 wraddr1 wraddr2 wraddr3 rdaddr0 rdaddr1 rdaddr2 rdaddr3 ESE370__Readaddr__Wraddr
XTristate@0 net@21 Last__write this__write ESE370__TristateBufferSized
VVPulse@3 net@208 gnd pulse (0 0.8 0ns 10ps 10ps 80ps 100ns) DC '0V' AC '0V' 0
XaddressL@0 wraddr3 wraddr2 wraddr1 wraddr0 clk willenq ESE370__addressLoop
XaddressL@1 rdaddr3 rdaddr2 rdaddr1 rdaddr0 clk willdq ESE370__addressLoop
Xand2@0 ptrflag net@43 Empty_next ESE370__and2
Xand2@1 ptrflag Last__write Full_next ESE370__and2
Xand2@2 ENQ andin willenq ESE370__and2
Xand2@3 DQ net@110 willdq ESE370__and2
Xand2@4 clk willenq net@287 ESE370__and2
Xbuffer@0 net@287 WRCtrl ESE370__buffer
Xinverter@1 Empty_next net@110 ESE370__inverter
Xinverter@2 Full_next andin ESE370__inverter
Xinverter@3 Last__write net@43 ESE370__inverter
Xnor2@0 willenq willdq net@21 ESE370__nor2
Xtristate@2 net@21 willenq this__write ESE370__tristate-buffer-enable-inverted
.ENDS ESE370__controlLogic

*** SUBCIRCUIT ESE370__tristate-inverter FROM CELL tristate-inverter{sch}
.SUBCKT ESE370__tristate-inverter En In out
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 out In net@13 gnd N L=0.022U W=0.022U
Mnmos@1 net@13 En gnd gnd N L=0.022U W=0.022U
Mpmos@0 net@0 In out vdd P L=0.022U W=0.022U
Mpmos@1 vdd net@28 net@0 vdd P L=0.022U W=0.022U
Xinverter@2 En net@28 ESE370__inverter
.ENDS ESE370__tristate-inverter

*** SUBCIRCUIT ESE370__dataDriver FROM CELL dataDriver{sch}
.SUBCKT ESE370__dataDriver bit0 bit1 bit2 bit3 d0 d0_ d1 d1_ d2 d2_ d3 d3_ En
** GLOBAL gnd
** GLOBAL vdd
Xtri-stat@0 En bit0 d0 ESE370__tri-state-buffer
Xtri-stat@1 En bit1 d1 ESE370__tri-state-buffer
Xtri-stat@2 En bit2 d2 ESE370__tri-state-buffer
Xtri-stat@3 En bit3 d3 ESE370__tri-state-buffer
Xtristate@4 En bit0 d0_ ESE370__tristate-inverter
Xtristate@5 En bit1 d1_ ESE370__tristate-inverter
Xtristate@6 En bit2 d2_ ESE370__tristate-inverter
Xtristate@7 En bit3 d3_ ESE370__tristate-inverter
.ENDS ESE370__dataDriver

*** SUBCIRCUIT ESE370__inputRegister FROM CELL inputRegister{sch}
.SUBCKT ESE370__inputRegister clk dequeue DQC enqueue EQC in0 in0C in1 in1C in2 in2C in3 in3C
** GLOBAL gnd
** GLOBAL vdd
X_4bitReg@0 clk in3 in2 in1 in0 in3C in2C in1C in0C ESE370__4bitReg
XPositive@0 clk enqueue EQC ESE370__PositiveRegister
XPositive@1 clk dequeue DQC ESE370__PositiveRegister
.ENDS ESE370__inputRegister

.global gnd vdd

*** TOP LEVEL CELL: SRAMtests{sch}
XSRAM@0 addr3 addr2 addr1 addr0 bl0 d3_ d2_ d1_ d0_ d3 d2 d1 d0 pc pcafter wl0 wl1 rw ESE370__SRAM
VVPWL@0 enqIn gnd pwl (0 0 2ns 0V 2ns 0.8V 6ns 0.8V 6ns 0V 8ns 0V) DC 0V AC 0V 0
VVPWL@1 DQIn gnd pwl (0 0 6ns 0V 6ns 0.8V 8ns 0.8V 8ns 0V 10ns 0V) DC 0V AC 0V 0
VVPulse@0 clk gnd pulse (0 0.8V 0ns 10ps 10ps 1ns 2ns) DC 0V AC 0V 0
VVPulse@1 pc gnd pulse (0.8V 0V 100ps 10ps 10ps 110ps 1ns) DC 0V AC 0V 0
VVPulse@2 in gnd pulse (0.8 0V 0ns 10ps 10ps 3.9ns 1s) DC 0V AC 0V 0
VV_Generi@0 vdd gnd DC 0.8 AC 0
XcontrolL@0 addr0 addr1 addr2 addr3 clk dq empty enq full rw ESE370__controlLogic
XdataDriv@0 in0 in1 in2 in3 d0 d0_ d1 d1_ d2 d2_ d3 d3_ rw ESE370__dataDriver
XinputReg@0 clk DQIn dq enqIn enq in in0 in in1 in in2 in in3 ESE370__inputRegister
.END
