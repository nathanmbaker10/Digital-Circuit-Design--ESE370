*** SPICE deck for cell SRAM{sch} from library ESE370
*** Created on Sun Nov 28, 2021 16:03:02
*** Last revised on Tue Nov 30, 2021 18:41:52
*** Written on Tue Nov 30, 2021 19:36:21 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF
* Model cards are described in this file:
.include '~/Desktop/Shared VM (Desktop)/ESE370/22nm_HP.pm'

*** SUBCIRCUIT ESE370__inverter FROM CELL inverter{sch}
.SUBCKT ESE370__inverter a not_a_
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 not_a_ a gnd gnd N L=0.022U W=0.022U
Mpmos@0 vdd a not_a_ vdd P L=0.022U W=0.022U
.ENDS ESE370__inverter

*** SUBCIRCUIT ESE370__buffer FROM CELL buffer{sch}
.SUBCKT ESE370__buffer a out
** GLOBAL gnd
** GLOBAL vdd
Xinverter@0 a net@1 ESE370__inverter
Xinverter@1 net@1 out ESE370__inverter
.ENDS ESE370__buffer

*** SUBCIRCUIT ESE370__ColumnChooser FROM CELL ColumnChooser{sch}
.SUBCKT ESE370__ColumnChooser C0 C1 In
** GLOBAL gnd
** GLOBAL vdd
Xbuffer@0 In C1 ESE370__buffer
Xinverter@0 In C0 ESE370__inverter
.ENDS ESE370__ColumnChooser

*** SUBCIRCUIT ESE370__tri-state-buffer FROM CELL tri-state-buffer{sch}
.SUBCKT ESE370__tri-state-buffer En In out
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 out En net@24 gnd N L=0.022U W=0.022U
Mnmos@1 net@24 net@3 gnd gnd N L=0.022U W=0.022U
Mpmos@0 net@1 net@14 out vdd P L=0.022U W=0.022U
Mpmos@1 vdd net@3 net@1 vdd P L=0.022U W=0.022U
Xinverter@1 In net@3 ESE370__inverter
Xinverter@2 En net@14 ESE370__inverter
.ENDS ESE370__tri-state-buffer

*** SUBCIRCUIT ESE370__TristateBufferSized FROM CELL TristateBufferSized{sch}
.SUBCKT ESE370__TristateBufferSized En In out
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 out En net@6 gnd N L=0.022U W=0.022U
Mnmos@1 net@6 net@10 gnd gnd N L=0.022U W=0.022U
Mpmos@0 net@1 net@17 out vdd P L=0.022U W=0.022U
Mpmos@1 vdd net@10 net@1 vdd P L=0.022U W=0.022U
Xinverter@0 In net@10 ESE370__inverter
Xinverter@1 En net@17 ESE370__inverter
.ENDS ESE370__TristateBufferSized

*** SUBCIRCUIT ESE370__tristateBufferEnableInvertedSized FROM CELL tristateBufferEnableInvertedSized{sch}
.SUBCKT ESE370__tristateBufferEnableInvertedSized En In out
** GLOBAL gnd
** GLOBAL vdd
XTristate@0 net@2 In out ESE370__TristateBufferSized
Xinverter@0 En net@2 ESE370__inverter
.ENDS ESE370__tristateBufferEnableInvertedSized

*** SUBCIRCUIT ESE370__ColumnDriver FROM CELL ColumnDriver{sch}
.SUBCKT ESE370__ColumnDriver b Cin d WR/_R
** GLOBAL gnd
** GLOBAL vdd
Xtri-stat@0 WR/_R d net@162 ESE370__tri-state-buffer
Xtri-stat@1 Cin net@162 b ESE370__tri-state-buffer
Xtri-stat@2 Cin b net@122 ESE370__tri-state-buffer
Xtristate@7 WR/_R net@122 d ESE370__tristateBufferEnableInvertedSized
.ENDS ESE370__ColumnDriver

*** SUBCIRCUIT ESE370__ColumnDecoderBus FROM CELL ColumnDecoderBus{sch}
.SUBCKT ESE370__ColumnDecoderBus BL_[7] BL_[6] BL_[5] BL_[4] BL_[3] BL_[2] BL_[1] BL_[0] BL[7] BL[6] BL[5] BL[4] BL[3] BL[2] BL[1] BL[0] Cin D_[3] D_[2] D_[1] D_[0] D[3] D[2] D[1] D[0] Wr/_R
** GLOBAL gnd
** GLOBAL vdd
XColumnCh@0 net@8 net@46 Cin ESE370__ColumnChooser
XColumnDr@0 BL[0] net@8 D[0] Wr/_R ESE370__ColumnDriver
XColumnDr@1 BL_[0] net@8 D_[0] Wr/_R ESE370__ColumnDriver
XColumnDr@4 BL[1] net@8 D[1] Wr/_R ESE370__ColumnDriver
XColumnDr@5 BL_[1] net@8 D_[1] Wr/_R ESE370__ColumnDriver
XColumnDr@6 BL[2] net@8 D[2] Wr/_R ESE370__ColumnDriver
XColumnDr@7 BL_[2] net@8 D_[2] Wr/_R ESE370__ColumnDriver
XColumnDr@8 BL[3] net@8 D[3] Wr/_R ESE370__ColumnDriver
XColumnDr@9 BL_[3] net@8 D_[3] Wr/_R ESE370__ColumnDriver
XColumnDr@10 BL[4] net@46 D[0] Wr/_R ESE370__ColumnDriver
XColumnDr@11 BL_[4] net@46 D_[0] Wr/_R ESE370__ColumnDriver
XColumnDr@12 BL[5] net@46 D[1] Wr/_R ESE370__ColumnDriver
XColumnDr@13 BL_[5] net@46 D_[1] Wr/_R ESE370__ColumnDriver
XColumnDr@14 BL[6] net@46 D[2] Wr/_R ESE370__ColumnDriver
XColumnDr@15 BL_[6] net@46 D_[2] Wr/_R ESE370__ColumnDriver
XColumnDr@16 BL[7] net@46 D[3] Wr/_R ESE370__ColumnDriver
XColumnDr@17 BL_[7] net@46 D_[3] Wr/_R ESE370__ColumnDriver
.ENDS ESE370__ColumnDecoderBus

*** SUBCIRCUIT ESE370__RAM_Cell FROM CELL RAM_Cell{sch}
.SUBCKT ESE370__RAM_Cell BL BL_ WL
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 net@0 WL BL gnd N L=0.022U W=0.044U
Mnmos@1 BL_ WL net@10 gnd N L=0.022U W=0.022U
Mnmos@2 net@10 net@0 gnd gnd N L=0.022U W=0.044U
Mnmos@3 net@0 net@10 gnd gnd N L=0.022U W=0.022U
Mpmos@0 vdd net@0 net@10 vdd P L=0.022U W=0.022U
Mpmos@1 vdd net@10 net@0 vdd P L=0.022U W=0.022U
.ENDS ESE370__RAM_Cell

*** SUBCIRCUIT ESE370__nand2 FROM CELL nand2{sch}
.SUBCKT ESE370__nand2 A B O
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 O A net@10 gnd N L=0.022U W=0.022U
Mnmos@1 net@10 B gnd gnd N L=0.022U W=0.022U
Mpmos@0 vdd A O vdd P L=0.022U W=0.022U
Mpmos@1 vdd B O vdd P L=0.022U W=0.022U
.ENDS ESE370__nand2

*** SUBCIRCUIT ESE370__and2 FROM CELL and2{sch}
.SUBCKT ESE370__and2 a b output
** GLOBAL gnd
** GLOBAL vdd
Xinverter@0 net@25 output ESE370__inverter
Xnand2@0 a b net@25 ESE370__nand2
.ENDS ESE370__and2

*** SUBCIRCUIT ESE370__RowDecoder FROM CELL RowDecoder{sch}
.SUBCKT ESE370__RowDecoder Addr[2] Addr[1] Addr[0] WL0 WL1 WL2 WL3 WL4 WL5 WL6 WL7 _PC
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 net@346 net@33 gnd gnd N L=0.022U W=0.022U
Mnmos@2 net@267 net@33 gnd gnd N L=0.022U W=0.022U
Mnmos@3 net@49 net@51 gnd gnd N L=0.022U W=0.022U
Mnmos@7 net@269 net@51 gnd gnd N L=0.022U W=0.022U
Mnmos@8 net@70 net@72 gnd gnd N L=0.022U W=0.022U
Mnmos@11 net@81 net@72 gnd gnd N L=0.022U W=0.022U
Mnmos@12 net@85 net@97 gnd gnd N L=0.022U W=0.022U
Mnmos@15 net@341 net@97 gnd gnd N L=0.022U W=0.022U
Mnmos@16 net@125 net@281 net@346 gnd N L=0.022U W=0.022U
Mnmos@17 net@130 Addr[0] net@267 gnd N L=0.022U W=0.022U
Mnmos@18 net@139 net@281 net@49 gnd N L=0.022U W=0.022U
Mnmos@19 net@145 Addr[0] net@269 gnd N L=0.022U W=0.022U
Mnmos@20 net@149 net@281 net@70 gnd N L=0.022U W=0.022U
Mnmos@21 net@153 Addr[0] net@81 gnd N L=0.022U W=0.022U
Mnmos@22 net@161 net@281 net@85 gnd N L=0.022U W=0.022U
Mnmos@23 net@94 Addr[0] net@341 gnd N L=0.022U W=0.022U
Mpmos@8 vdd _PC net@125 vdd P L=0.022U W=0.044U
Mpmos@9 vdd _PC net@130 vdd P L=0.022U W=0.044U
Mpmos@10 vdd _PC net@139 vdd P L=0.022U W=0.044U
Mpmos@11 vdd _PC net@145 vdd P L=0.022U W=0.044U
Mpmos@12 vdd _PC net@149 vdd P L=0.022U W=0.044U
Mpmos@13 vdd _PC net@153 vdd P L=0.022U W=0.044U
Mpmos@14 vdd _PC net@161 vdd P L=0.022U W=0.044U
Mpmos@15 vdd _PC net@94 vdd P L=0.022U W=0.044U
Xand2@0 Addr[1] Addr[2] net@97 ESE370__and2
Xand2@1 net@10 Addr[2] net@51 ESE370__and2
Xand2@2 Addr[1] net@9 net@72 ESE370__and2
Xand2@3 net@8 net@7 net@33 ESE370__and2
Xinverter@1 Addr[2] net@7 ESE370__inverter
Xinverter@2 Addr[1] net@8 ESE370__inverter
Xinverter@3 Addr[2] net@9 ESE370__inverter
Xinverter@4 Addr[1] net@10 ESE370__inverter
Xinverter@6 net@125 WL0 ESE370__inverter
Xinverter@7 net@130 WL1 ESE370__inverter
Xinverter@8 net@139 WL2 ESE370__inverter
Xinverter@9 net@145 WL3 ESE370__inverter
Xinverter@10 net@149 WL4 ESE370__inverter
Xinverter@11 net@153 WL5 ESE370__inverter
Xinverter@12 net@161 WL6 ESE370__inverter
Xinverter@13 net@94 WL7 ESE370__inverter
Xinverter@14 Addr[0] net@281 ESE370__inverter
.ENDS ESE370__RowDecoder

*** SUBCIRCUIT ESE370__bitLineConditioning FROM CELL bitLineConditioning{sch}
.SUBCKT ESE370__bitLineConditioning BL BL_ CLK
** GLOBAL vdd
Mpmos@0 vdd CLK BL_ vdd P L=0.022U W=0.022U
Mpmos@2 vdd CLK BL vdd P L=0.022U W=0.022U
.ENDS ESE370__bitLineConditioning

*** SUBCIRCUIT ESE370__tristate-inverter FROM CELL tristate-inverter{sch}
.SUBCKT ESE370__tristate-inverter En In out
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 out In net@13 gnd N L=0.022U W=0.022U
Mnmos@1 net@13 En gnd gnd N L=0.022U W=0.022U
Mpmos@0 net@0 In out vdd P L=0.022U W=0.022U
Mpmos@1 vdd net@28 net@0 vdd P L=0.022U W=0.022U
Xinverter@2 En net@28 ESE370__inverter
.ENDS ESE370__tristate-inverter

*** SUBCIRCUIT ESE370__tristate-buffer-enable-inverted FROM CELL tristate-buffer-enable-inverted{sch}
.SUBCKT ESE370__tristate-buffer-enable-inverted en in out
** GLOBAL gnd
** GLOBAL vdd
Xinverter@0 en net@2 ESE370__inverter
Xtri-stat@0 net@2 in out ESE370__tri-state-buffer
.ENDS ESE370__tristate-buffer-enable-inverted

.global gnd vdd

*** TOP LEVEL CELL: SRAM{sch}
XColumnDe@0 net@161 net@147 net@133 net@119 bl_4 bl_3 bl_2 bl_ net@154 net@140 net@126 net@112 bl4 bl3 bl2 bl gnd gnd gnd gnd Q_ gnd gnd gnd Q RW ESE370__ColumnDecoderBus
XRAM_Cell@0 bl bl_ wl0 ESE370__RAM_Cell
XRAM_Cell@1 bl2 bl_2 wl0 ESE370__RAM_Cell
XRAM_Cell@2 bl3 bl_3 wl0 ESE370__RAM_Cell
XRAM_Cell@3 bl4 bl_4 wl0 ESE370__RAM_Cell
XRAM_Cell@8 net@112 net@119 wl0 ESE370__RAM_Cell
XRAM_Cell@9 net@126 net@133 wl0 ESE370__RAM_Cell
XRAM_Cell@10 net@140 net@147 wl0 ESE370__RAM_Cell
XRAM_Cell@11 net@154 net@161 wl0 ESE370__RAM_Cell
XRAM_Cell@12 bl bl_ wl1 ESE370__RAM_Cell
XRAM_Cell@13 bl2 bl_2 wl1 ESE370__RAM_Cell
XRAM_Cell@14 bl3 bl_3 wl1 ESE370__RAM_Cell
XRAM_Cell@15 bl4 bl_4 wl1 ESE370__RAM_Cell
XRAM_Cell@16 net@112 net@119 wl1 ESE370__RAM_Cell
XRAM_Cell@17 net@126 net@133 wl1 ESE370__RAM_Cell
XRAM_Cell@18 net@140 net@147 wl1 ESE370__RAM_Cell
XRAM_Cell@19 net@154 net@161 wl1 ESE370__RAM_Cell
XRAM_Cell@20 bl bl_ wl2 ESE370__RAM_Cell
XRAM_Cell@21 bl2 bl_2 wl2 ESE370__RAM_Cell
XRAM_Cell@22 bl3 bl_3 wl2 ESE370__RAM_Cell
XRAM_Cell@23 bl4 bl_4 wl2 ESE370__RAM_Cell
XRAM_Cell@24 net@112 net@119 wl2 ESE370__RAM_Cell
XRAM_Cell@25 net@126 net@133 wl2 ESE370__RAM_Cell
XRAM_Cell@26 net@140 net@147 wl2 ESE370__RAM_Cell
XRAM_Cell@27 net@154 net@161 wl2 ESE370__RAM_Cell
XRAM_Cell@28 bl bl_ wl3 ESE370__RAM_Cell
XRAM_Cell@29 bl2 bl_2 wl3 ESE370__RAM_Cell
XRAM_Cell@30 bl3 bl_3 wl3 ESE370__RAM_Cell
XRAM_Cell@31 bl4 bl_4 wl3 ESE370__RAM_Cell
XRAM_Cell@32 net@112 net@119 wl3 ESE370__RAM_Cell
XRAM_Cell@33 net@126 net@133 wl3 ESE370__RAM_Cell
XRAM_Cell@34 net@140 net@147 wl3 ESE370__RAM_Cell
XRAM_Cell@35 net@154 net@161 wl3 ESE370__RAM_Cell
XRAM_Cell@36 bl bl_ wl4 ESE370__RAM_Cell
XRAM_Cell@37 bl2 bl_2 wl4 ESE370__RAM_Cell
XRAM_Cell@38 bl3 bl_3 wl4 ESE370__RAM_Cell
XRAM_Cell@39 bl4 bl_4 wl4 ESE370__RAM_Cell
XRAM_Cell@40 net@112 net@119 wl4 ESE370__RAM_Cell
XRAM_Cell@41 net@126 net@133 wl4 ESE370__RAM_Cell
XRAM_Cell@42 net@140 net@147 wl4 ESE370__RAM_Cell
XRAM_Cell@43 net@154 net@161 wl4 ESE370__RAM_Cell
XRAM_Cell@44 bl bl_ wl5 ESE370__RAM_Cell
XRAM_Cell@45 bl2 bl_2 wl5 ESE370__RAM_Cell
XRAM_Cell@46 bl3 bl_3 wl5 ESE370__RAM_Cell
XRAM_Cell@47 bl4 bl_4 wl5 ESE370__RAM_Cell
XRAM_Cell@48 net@112 net@119 wl5 ESE370__RAM_Cell
XRAM_Cell@49 net@126 net@133 wl5 ESE370__RAM_Cell
XRAM_Cell@50 net@140 net@147 wl5 ESE370__RAM_Cell
XRAM_Cell@51 net@154 net@161 wl5 ESE370__RAM_Cell
XRAM_Cell@52 bl bl_ wl6 ESE370__RAM_Cell
XRAM_Cell@53 bl2 bl_2 wl6 ESE370__RAM_Cell
XRAM_Cell@54 bl3 bl_3 wl6 ESE370__RAM_Cell
XRAM_Cell@55 bl4 bl_4 wl6 ESE370__RAM_Cell
XRAM_Cell@56 net@112 net@119 wl6 ESE370__RAM_Cell
XRAM_Cell@57 net@126 net@133 wl6 ESE370__RAM_Cell
XRAM_Cell@58 net@140 net@147 wl6 ESE370__RAM_Cell
XRAM_Cell@59 net@154 net@161 wl6 ESE370__RAM_Cell
XRAM_Cell@60 bl bl_ wl7 ESE370__RAM_Cell
XRAM_Cell@61 bl2 bl_2 wl7 ESE370__RAM_Cell
XRAM_Cell@62 bl3 bl_3 wl7 ESE370__RAM_Cell
XRAM_Cell@63 bl4 bl_4 wl7 ESE370__RAM_Cell
XRAM_Cell@64 net@112 net@119 wl7 ESE370__RAM_Cell
XRAM_Cell@65 net@126 net@133 wl7 ESE370__RAM_Cell
XRAM_Cell@66 net@140 net@147 wl7 ESE370__RAM_Cell
XRAM_Cell@67 net@154 net@161 wl7 ESE370__RAM_Cell
XRowDecod@4 gnd gnd gnd wl0 wl1 wl2 wl3 wl4 wl5 wl6 wl7 pcbefore ESE370__RowDecoder
VVPWL@0 net@302 gnd pwl (0ns 0.8 1ns 0.8 1ns 0 2.667ns 0 2.667ns 0.8) DC 0V AC 0V 0
VVPulse@0 pcbefore gnd pulse (0.8V 0V 20ps 10ps 10ps 110ps 333ps) DC 0V AC 0V 0
VVPulse@1 RW gnd pulse (0V 0.8V 0ps 10ps 10ps 333ps 1ns) DC 0V AC 0V 0
VV_Generi@0 vdd gnd DC 0.8 AC 0
XbitLineC@0 bl bl_ pcafter ESE370__bitLineConditioning
XbitLineC@1 bl2 bl_2 pcafter ESE370__bitLineConditioning
XbitLineC@2 bl3 bl_3 pcafter ESE370__bitLineConditioning
XbitLineC@3 bl4 bl_4 pcafter ESE370__bitLineConditioning
XbitLineC@4 net@112 net@119 pcafter ESE370__bitLineConditioning
XbitLineC@5 net@126 net@133 pcafter ESE370__bitLineConditioning
XbitLineC@7 net@140 net@147 pcafter ESE370__bitLineConditioning
XbitLineC@8 net@154 net@161 pcafter ESE370__bitLineConditioning
Xtri-stat@0 RW net@302 Q ESE370__tri-state-buffer
Xtristate@0 RW net@302 Q_ ESE370__tristate-inverter
Xtristate@1 RW pcbefore pcafter ESE370__tristate-buffer-enable-inverted
.END
