*** SPICE deck for cell HW6Q2{sch} from library ESE370
*** Created on Wed Nov 10, 2021 22:37:51
*** Last revised on Thu Nov 11, 2021 21:18:25
*** Written on Thu Nov 11, 2021 21:21:42 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF
* Model cards are described in this file:
.include '~/Desktop/Shared VM (Desktop)/ESE370/22nm_HP.pm'

*** SUBCIRCUIT ESE370__inverter FROM CELL inverter{sch}
.SUBCKT ESE370__inverter a not_a_
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 not_a_ a gnd gnd N L=0.022U W=0.022U
Mpmos@0 vdd a not_a_ vdd P L=0.022U W=0.022U
.ENDS ESE370__inverter

*** SUBCIRCUIT ESE370__nand2 FROM CELL nand2{sch}
.SUBCKT ESE370__nand2 A B O
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 O A net@10 gnd N L=0.022U W=0.022U
Mnmos@1 net@10 B gnd gnd N L=0.022U W=0.022U
Mpmos@0 vdd A O vdd P L=0.022U W=0.022U
Mpmos@1 vdd B O vdd P L=0.022U W=0.022U
.ENDS ESE370__nand2

*** SUBCIRCUIT ESE370__3nandlatch FROM CELL 3nandlatch{sch}
.SUBCKT ESE370__3nandlatch clock in out
** GLOBAL gnd
** GLOBAL vdd
Xinverter@0 clock net@6 ESE370__inverter
Xnand2@0 in clock net@8 ESE370__nand2
Xnand2@1 net@6 out net@10 ESE370__nand2
Xnand2@2 net@8 net@10 out ESE370__nand2
.ENDS ESE370__3nandlatch

.global gnd vdd

*** TOP LEVEL CELL: HW6Q2{sch}
X_3nandlat@0 vdd net@7 net@9 ESE370__3nandlatch
X_3nandlat@1 _3nandlat@1_clock net@9 _3nandlat@1_out ESE370__3nandlatch
VVPulse@1 net@7 gnd pulse (0 0.8V 0ns 10ps 10ps 1.5ns 3ns) DC '0V' AC '0V' 0
VV_Generi@0 vdd gnd 'DC 0.8 AC 0'
.END
